module juego(input logic up,
input logic down,
input logic right,
input logic left,
input logic play,
input logic reset,
input logic clk,
output reg[15:0] PairsCards,
output reg[15:0] OpenCards,
output reg[1:0] win,
output logic timeOut);



endmodule